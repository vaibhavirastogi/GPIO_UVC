`include "uvm_macros.svh"
import uvm_pkg::*;
`include "def.sv"  
`include "gpio_seq_item.sv"
`include "gpio_seq_item_ext.sv"
`include "gpio_sequencer.sv"
`include "gpio_sequence.sv"
`include "gpio_driver.sv"
`include "gpio_trans_item.sv"
`include "gpio_monitor.sv"
`include "gpio_agent.sv"
`include "gpio_env.sv"
`include "agent_config.sv"
`include "agent_config_ext.sv"
`include "gpio_test.sv"
