`define MAX_SYNCINPUT 16
`define MAX_SYNCOUTPUT 16
`define MAX_ASYNCINPUT 16
`define MAX_ASYNCOUTPUT 16
`define MAX_SYNCOP 16
`define MAX_ASYNCOP 16
`define NO_TRANSCATION 50
